//ディスプレイ固有の設定値とか保管

parameter VPERIOD  = 10'd112;
parameter VFRONT   = 10'd16;
parameter VWIDTH   = 10'd96;
parameter VBACK    = 10'd0;

parameter HPERIOD  = 10'd507;
parameter HFRONT   = 10'd107;
parameter HWIDTH   = 10'd400;
parameter HBACK    = 10'd0;
